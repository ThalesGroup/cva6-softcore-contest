// Copyright 2018 ETH Zurich and University of Bologna.
// Copyright and related rights are licensed under the Solderpad Hardware
// License, Version 0.51 (the "License"); you may not use this file except in
// compliance with the License.  You may obtain a copy of the License at
// http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
// or agreed to in writing, software, hardware and materials distributed under
// this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
// CONDITIONS OF ANY KIND, either express or implied. See the License for the
// specific language governing permissions and limitations under the License.

// Xilinx Peripherals

`include "axi/assign.svh"
`include "axi/typedef.svh"
`include "register_interface/assign.svh"
`include "register_interface/typedef.svh"

module ariane_peripherals #(
  parameter int AxiAddrWidth = -1,
  parameter int AxiDataWidth = -1,
  parameter int AxiIdWidth   = -1,
  parameter int AxiUserWidth = 1,
  parameter bit InclUART     = 1,
  parameter bit InclSPI      = 0,
  parameter bit InclEthernet = 0,
  parameter bit InclGPIO     = 0,
  parameter bit InclTimer    = 1,
  //VGA
  parameter int unsigned RedWidth     = 5,
  parameter int unsigned GreenWidth   = 6,
  parameter int unsigned BlueWidth    = 5,
  parameter int unsigned HCountWidth  = 32,
  parameter int unsigned VCountWidth  = 32
) (
  input  logic       clk_i,           // Clock
  input  logic       clk_200MHz_i,
  input  logic       clk_vga_i,
  input  logic       rst_ni,          // Asynchronous reset active low
  AXI_BUS.Slave      plic,
  AXI_BUS.Slave      uart,
  AXI_BUS.Slave      spi,
  AXI_BUS.Slave      gpio,
  AXI_BUS.Slave      ethernet,
  AXI_BUS.Slave      timer,
  AXI_BUS.Slave      vga, 
  AXI_BUS.Master     mvga,
  output logic [1:0] irq_o,
  // UART
  input  logic       rx_i,
  output logic       tx_o,
  // Ethernet
  input  logic       eth_clk_i,
  input  wire        eth_rxck,
  input  wire        eth_rxctl,
  input  wire [3:0]  eth_rxd,
  output wire        eth_txck,
  output wire        eth_txctl,
  output wire [3:0]  eth_txd,
  output wire        eth_rst_n,
  input  logic       phy_tx_clk_i,    // 125 MHz Clock
  // MDIO Interface
  inout  wire        eth_mdio,
  output logic       eth_mdc,
  // SPI
  output logic       spi_clk_o,
  output logic       spi_mosi,
  input  logic       spi_miso,
  output logic       spi_ss,
  // SD Card
  input  logic       sd_clk_i,
  output logic [7:0] leds_o,
  input  logic [7:0] dip_switches_i,
  // VGA
  output logic                  hsync,
  output logic                  vsync,
  output logic [RedWidth-1:0]   red,
  output logic [GreenWidth-1:0] green,
  output logic [BlueWidth-1:0]  blue
);

  // ---------------
  // 1. PLIC
  // ---------------
  logic [ariane_soc::NumSources-1:0] irq_sources;

  // Unused interrupt sources
  assign irq_sources[ariane_soc::NumSources-1:8] = '0;

  REG_BUS #(
    .ADDR_WIDTH ( 32 ),
    .DATA_WIDTH ( 32 )
  ) reg_bus (clk_i);

  logic         plic_penable;
  logic         plic_pwrite;
  logic [31:0]  plic_paddr;
  logic         plic_psel;
  logic [31:0]  plic_pwdata;
  logic [31:0]  plic_prdata;
  logic         plic_pready;
  logic         plic_pslverr;

  axi2apb_64_32 #(
    .AXI4_ADDRESS_WIDTH ( AxiAddrWidth  ),
    .AXI4_RDATA_WIDTH   ( AxiDataWidth  ),
    .AXI4_WDATA_WIDTH   ( AxiDataWidth  ),
    .AXI4_ID_WIDTH      ( AxiIdWidth    ),
    .AXI4_USER_WIDTH    ( AxiUserWidth  ),
    .BUFF_DEPTH_SLAVE   ( 2             ),
    .APB_ADDR_WIDTH     ( 32            )
  ) i_axi2apb_64_32_plic (
    .ACLK      ( clk_i          ),
    .ARESETn   ( rst_ni         ),
    .test_en_i ( 1'b0           ),
    .AWID_i    ( plic.aw_id     ),
    .AWADDR_i  ( plic.aw_addr   ),
    .AWLEN_i   ( plic.aw_len    ),
    .AWSIZE_i  ( plic.aw_size   ),
    .AWBURST_i ( plic.aw_burst  ),
    .AWLOCK_i  ( plic.aw_lock   ),
    .AWCACHE_i ( plic.aw_cache  ),
    .AWPROT_i  ( plic.aw_prot   ),
    .AWREGION_i( plic.aw_region ),
    .AWUSER_i  ( plic.aw_user   ),
    .AWQOS_i   ( plic.aw_qos    ),
    .AWVALID_i ( plic.aw_valid  ),
    .AWREADY_o ( plic.aw_ready  ),
    .WDATA_i   ( plic.w_data    ),
    .WSTRB_i   ( plic.w_strb    ),
    .WLAST_i   ( plic.w_last    ),
    .WUSER_i   ( plic.w_user    ),
    .WVALID_i  ( plic.w_valid   ),
    .WREADY_o  ( plic.w_ready   ),
    .BID_o     ( plic.b_id      ),
    .BRESP_o   ( plic.b_resp    ),
    .BVALID_o  ( plic.b_valid   ),
    .BUSER_o   ( plic.b_user    ),
    .BREADY_i  ( plic.b_ready   ),
    .ARID_i    ( plic.ar_id     ),
    .ARADDR_i  ( plic.ar_addr   ),
    .ARLEN_i   ( plic.ar_len    ),
    .ARSIZE_i  ( plic.ar_size   ),
    .ARBURST_i ( plic.ar_burst  ),
    .ARLOCK_i  ( plic.ar_lock   ),
    .ARCACHE_i ( plic.ar_cache  ),
    .ARPROT_i  ( plic.ar_prot   ),
    .ARREGION_i( plic.ar_region ),
    .ARUSER_i  ( plic.ar_user   ),
    .ARQOS_i   ( plic.ar_qos    ),
    .ARVALID_i ( plic.ar_valid  ),
    .ARREADY_o ( plic.ar_ready  ),
    .RID_o     ( plic.r_id      ),
    .RDATA_o   ( plic.r_data    ),
    .RRESP_o   ( plic.r_resp    ),
    .RLAST_o   ( plic.r_last    ),
    .RUSER_o   ( plic.r_user    ),
    .RVALID_o  ( plic.r_valid   ),
    .RREADY_i  ( plic.r_ready   ),
    .PENABLE   ( plic_penable   ),
    .PWRITE    ( plic_pwrite    ),
    .PADDR     ( plic_paddr     ),
    .PSEL      ( plic_psel      ),
    .PWDATA    ( plic_pwdata    ),
    .PRDATA    ( plic_prdata    ),
    .PREADY    ( plic_pready    ),
    .PSLVERR   ( plic_pslverr   )
  );

  apb_to_reg i_apb_to_reg (
    .clk_i     ( clk_i        ),
    .rst_ni    ( rst_ni       ),
    .penable_i ( plic_penable ),
    .pwrite_i  ( plic_pwrite  ),
    .paddr_i   ( plic_paddr   ),
    .psel_i    ( plic_psel    ),
    .pwdata_i  ( plic_pwdata  ),
    .prdata_o  ( plic_prdata  ),
    .pready_o  ( plic_pready  ),
    .pslverr_o ( plic_pslverr ),
    .reg_o     ( reg_bus      )
  );

  // define reg type according to REG_BUS above
  `REG_BUS_TYPEDEF_ALL(plic, logic[31:0], logic[31:0], logic[3:0])
  plic_req_t plic_req;
  plic_rsp_t plic_rsp;

  // assign REG_BUS.out to (req_t, rsp_t) pair
  `REG_BUS_ASSIGN_TO_REQ(plic_req, reg_bus)
  `REG_BUS_ASSIGN_FROM_RSP(reg_bus, plic_rsp)

  plic_top #(
    .N_SOURCE    ( ariane_soc::NumSources  ),
    .N_TARGET    ( ariane_soc::NumTargets  ),
    .MAX_PRIO    ( ariane_soc::MaxPriority ),
    .reg_req_t   ( plic_req_t              ),
    .reg_rsp_t   ( plic_rsp_t              )
  ) i_plic (
    .clk_i,
    .rst_ni,
    .req_i         ( plic_req    ),
    .resp_o        ( plic_rsp    ),
    .le_i          ( '0          ), // 0:level 1:edge
    .irq_sources_i ( irq_sources ),
    .eip_targets_o ( irq_o       )
  );

  // ---------------
  // 2. UART
  // ---------------
  logic         uart_penable;
  logic         uart_pwrite;
  logic [31:0]  uart_paddr;
  logic         uart_psel;
  logic [31:0]  uart_pwdata;
  logic [31:0]  uart_prdata;
  logic         uart_pready;
  logic         uart_pslverr;

  axi2apb_64_32 #(
    .AXI4_ADDRESS_WIDTH ( AxiAddrWidth ),
    .AXI4_RDATA_WIDTH   ( AxiDataWidth ),
    .AXI4_WDATA_WIDTH   ( AxiDataWidth ),
    .AXI4_ID_WIDTH      ( AxiIdWidth   ),
    .AXI4_USER_WIDTH    ( AxiUserWidth ),
    .BUFF_DEPTH_SLAVE   ( 2            ),
    .APB_ADDR_WIDTH     ( 32           )
  ) i_axi2apb_64_32_uart (
    .ACLK      ( clk_i          ),
    .ARESETn   ( rst_ni         ),
    .test_en_i ( 1'b0           ),
    .AWID_i    ( uart.aw_id     ),
    .AWADDR_i  ( uart.aw_addr   ),
    .AWLEN_i   ( uart.aw_len    ),
    .AWSIZE_i  ( uart.aw_size   ),
    .AWBURST_i ( uart.aw_burst  ),
    .AWLOCK_i  ( uart.aw_lock   ),
    .AWCACHE_i ( uart.aw_cache  ),
    .AWPROT_i  ( uart.aw_prot   ),
    .AWREGION_i( uart.aw_region ),
    .AWUSER_i  ( uart.aw_user   ),
    .AWQOS_i   ( uart.aw_qos    ),
    .AWVALID_i ( uart.aw_valid  ),
    .AWREADY_o ( uart.aw_ready  ),
    .WDATA_i   ( uart.w_data    ),
    .WSTRB_i   ( uart.w_strb    ),
    .WLAST_i   ( uart.w_last    ),
    .WUSER_i   ( uart.w_user    ),
    .WVALID_i  ( uart.w_valid   ),
    .WREADY_o  ( uart.w_ready   ),
    .BID_o     ( uart.b_id      ),
    .BRESP_o   ( uart.b_resp    ),
    .BVALID_o  ( uart.b_valid   ),
    .BUSER_o   ( uart.b_user    ),
    .BREADY_i  ( uart.b_ready   ),
    .ARID_i    ( uart.ar_id     ),
    .ARADDR_i  ( uart.ar_addr   ),
    .ARLEN_i   ( uart.ar_len    ),
    .ARSIZE_i  ( uart.ar_size   ),
    .ARBURST_i ( uart.ar_burst  ),
    .ARLOCK_i  ( uart.ar_lock   ),
    .ARCACHE_i ( uart.ar_cache  ),
    .ARPROT_i  ( uart.ar_prot   ),
    .ARREGION_i( uart.ar_region ),
    .ARUSER_i  ( uart.ar_user   ),
    .ARQOS_i   ( uart.ar_qos    ),
    .ARVALID_i ( uart.ar_valid  ),
    .ARREADY_o ( uart.ar_ready  ),
    .RID_o     ( uart.r_id      ),
    .RDATA_o   ( uart.r_data    ),
    .RRESP_o   ( uart.r_resp    ),
    .RLAST_o   ( uart.r_last    ),
    .RUSER_o   ( uart.r_user    ),
    .RVALID_o  ( uart.r_valid   ),
    .RREADY_i  ( uart.r_ready   ),
    .PENABLE   ( uart_penable   ),
    .PWRITE    ( uart_pwrite    ),
    .PADDR     ( uart_paddr     ),
    .PSEL      ( uart_psel      ),
    .PWDATA    ( uart_pwdata    ),
    .PRDATA    ( uart_prdata    ),
    .PREADY    ( uart_pready    ),
    .PSLVERR   ( uart_pslverr   )
  );

  if (InclUART) begin : gen_uart
    apb_uart i_apb_uart (
      .CLK     ( clk_i           ),
      .RSTN    ( rst_ni          ),
      .PSEL    ( uart_psel       ),
      .PENABLE ( uart_penable    ),
      .PWRITE  ( uart_pwrite     ),
      .PADDR   ( uart_paddr[4:2] ),
      .PWDATA  ( uart_pwdata     ),
      .PRDATA  ( uart_prdata     ),
      .PREADY  ( uart_pready     ),
      .PSLVERR ( uart_pslverr    ),
      .INT     ( irq_sources[0]  ),
      .OUT1N   (                 ), // keep open
      .OUT2N   (                 ), // keep open
      .RTSN    (                 ), // no flow control
      .DTRN    (                 ), // no flow control
      .CTSN    ( 1'b0            ),
      .DSRN    ( 1'b0            ),
      .DCDN    ( 1'b0            ),
      .RIN     ( 1'b0            ),
      .SIN     ( rx_i            ),
      .SOUT    ( tx_o            )
    );
  end else begin
    /* pragma translate_off */
    `ifndef VERILATOR
    mock_uart i_mock_uart (
      .clk_i     ( clk_i        ),
      .rst_ni    ( rst_ni       ),
      .penable_i ( uart_penable ),
      .pwrite_i  ( uart_pwrite  ),
      .paddr_i   ( uart_paddr   ),
      .psel_i    ( uart_psel    ),
      .pwdata_i  ( uart_pwdata  ),
      .prdata_o  ( uart_prdata  ),
      .pready_o  ( uart_pready  ),
      .pslverr_o ( uart_pslverr )
    );
    `endif
    /* pragma translate_on */
  end

  // ---------------
  // 3. SPI
  // ---------------
  assign spi.b_user = 1'b0;
  assign spi.r_user = 1'b0;

  if (InclSPI) begin : gen_spi
    logic [31:0] s_axi_spi_awaddr;
    logic [7:0]  s_axi_spi_awlen;
    logic [2:0]  s_axi_spi_awsize;
    logic [1:0]  s_axi_spi_awburst;
    logic [0:0]  s_axi_spi_awlock;
    logic [3:0]  s_axi_spi_awcache;
    logic [2:0]  s_axi_spi_awprot;
    logic [3:0]  s_axi_spi_awregion;
    logic [3:0]  s_axi_spi_awqos;
    logic        s_axi_spi_awvalid;
    logic        s_axi_spi_awready;
    logic [31:0] s_axi_spi_wdata;
    logic [3:0]  s_axi_spi_wstrb;
    logic        s_axi_spi_wlast;
    logic        s_axi_spi_wvalid;
    logic        s_axi_spi_wready;
    logic [1:0]  s_axi_spi_bresp;
    logic        s_axi_spi_bvalid;
    logic        s_axi_spi_bready;
    logic [31:0] s_axi_spi_araddr;
    logic [7:0]  s_axi_spi_arlen;
    logic [2:0]  s_axi_spi_arsize;
    logic [1:0]  s_axi_spi_arburst;
    logic [0:0]  s_axi_spi_arlock;
    logic [3:0]  s_axi_spi_arcache;
    logic [2:0]  s_axi_spi_arprot;
    logic [3:0]  s_axi_spi_arregion;
    logic [3:0]  s_axi_spi_arqos;
    logic        s_axi_spi_arvalid;
    logic        s_axi_spi_arready;
    logic [31:0] s_axi_spi_rdata;
    logic [1:0]  s_axi_spi_rresp;
    logic        s_axi_spi_rlast;
    logic        s_axi_spi_rvalid;
    logic        s_axi_spi_rready;

    xlnx_axi_dwidth_converter i_xlnx_axi_dwidth_converter_spi (
      .s_axi_aclk     ( clk_i              ),
      .s_axi_aresetn  ( rst_ni             ),
      .s_axi_awid     ( spi.aw_id          ),
      .s_axi_awaddr   ( spi.aw_addr[31:0]  ),
      .s_axi_awlen    ( spi.aw_len         ),
      .s_axi_awsize   ( spi.aw_size        ),
      .s_axi_awburst  ( spi.aw_burst       ),
      .s_axi_awlock   ( spi.aw_lock        ),
      .s_axi_awcache  ( spi.aw_cache       ),
      .s_axi_awprot   ( spi.aw_prot        ),
      .s_axi_awregion ( spi.aw_region      ),
      .s_axi_awqos    ( spi.aw_qos         ),
      .s_axi_awvalid  ( spi.aw_valid       ),
      .s_axi_awready  ( spi.aw_ready       ),
      .s_axi_wdata    ( spi.w_data         ),
      .s_axi_wstrb    ( spi.w_strb         ),
      .s_axi_wlast    ( spi.w_last         ),
      .s_axi_wvalid   ( spi.w_valid        ),
      .s_axi_wready   ( spi.w_ready        ),
      .s_axi_bid      ( spi.b_id           ),
      .s_axi_bresp    ( spi.b_resp         ),
      .s_axi_bvalid   ( spi.b_valid        ),
      .s_axi_bready   ( spi.b_ready        ),
      .s_axi_arid     ( spi.ar_id          ),
      .s_axi_araddr   ( spi.ar_addr[31:0]  ),
      .s_axi_arlen    ( spi.ar_len         ),
      .s_axi_arsize   ( spi.ar_size        ),
      .s_axi_arburst  ( spi.ar_burst       ),
      .s_axi_arlock   ( spi.ar_lock        ),
      .s_axi_arcache  ( spi.ar_cache       ),
      .s_axi_arprot   ( spi.ar_prot        ),
      .s_axi_arregion ( spi.ar_region      ),
      .s_axi_arqos    ( spi.ar_qos         ),
      .s_axi_arvalid  ( spi.ar_valid       ),
      .s_axi_arready  ( spi.ar_ready       ),
      .s_axi_rid      ( spi.r_id           ),
      .s_axi_rdata    ( spi.r_data         ),
      .s_axi_rresp    ( spi.r_resp         ),
      .s_axi_rlast    ( spi.r_last         ),
      .s_axi_rvalid   ( spi.r_valid        ),
      .s_axi_rready   ( spi.r_ready        ),

      .m_axi_awaddr   ( s_axi_spi_awaddr   ),
      .m_axi_awlen    ( s_axi_spi_awlen    ),
      .m_axi_awsize   ( s_axi_spi_awsize   ),
      .m_axi_awburst  ( s_axi_spi_awburst  ),
      .m_axi_awlock   ( s_axi_spi_awlock   ),
      .m_axi_awcache  ( s_axi_spi_awcache  ),
      .m_axi_awprot   ( s_axi_spi_awprot   ),
      .m_axi_awregion ( s_axi_spi_awregion ),
      .m_axi_awqos    ( s_axi_spi_awqos    ),
      .m_axi_awvalid  ( s_axi_spi_awvalid  ),
      .m_axi_awready  ( s_axi_spi_awready  ),
      .m_axi_wdata    ( s_axi_spi_wdata    ),
      .m_axi_wstrb    ( s_axi_spi_wstrb    ),
      .m_axi_wlast    ( s_axi_spi_wlast    ),
      .m_axi_wvalid   ( s_axi_spi_wvalid   ),
      .m_axi_wready   ( s_axi_spi_wready   ),
      .m_axi_bresp    ( s_axi_spi_bresp    ),
      .m_axi_bvalid   ( s_axi_spi_bvalid   ),
      .m_axi_bready   ( s_axi_spi_bready   ),
      .m_axi_araddr   ( s_axi_spi_araddr   ),
      .m_axi_arlen    ( s_axi_spi_arlen    ),
      .m_axi_arsize   ( s_axi_spi_arsize   ),
      .m_axi_arburst  ( s_axi_spi_arburst  ),
      .m_axi_arlock   ( s_axi_spi_arlock   ),
      .m_axi_arcache  ( s_axi_spi_arcache  ),
      .m_axi_arprot   ( s_axi_spi_arprot   ),
      .m_axi_arregion ( s_axi_spi_arregion ),
      .m_axi_arqos    ( s_axi_spi_arqos    ),
      .m_axi_arvalid  ( s_axi_spi_arvalid  ),
      .m_axi_arready  ( s_axi_spi_arready  ),
      .m_axi_rdata    ( s_axi_spi_rdata    ),
      .m_axi_rresp    ( s_axi_spi_rresp    ),
      .m_axi_rlast    ( s_axi_spi_rlast    ),
      .m_axi_rvalid   ( s_axi_spi_rvalid   ),
      .m_axi_rready   ( s_axi_spi_rready   )
    );

    xlnx_axi_quad_spi i_xlnx_axi_quad_spi (
      .ext_spi_clk    ( clk_i                  ),
      .s_axi4_aclk    ( clk_i                  ),
      .s_axi4_aresetn ( rst_ni                 ),
      .s_axi4_awaddr  ( s_axi_spi_awaddr[23:0] ),
      .s_axi4_awlen   ( s_axi_spi_awlen        ),
      .s_axi4_awsize  ( s_axi_spi_awsize       ),
      .s_axi4_awburst ( s_axi_spi_awburst      ),
      .s_axi4_awlock  ( s_axi_spi_awlock       ),
      .s_axi4_awcache ( s_axi_spi_awcache      ),
      .s_axi4_awprot  ( s_axi_spi_awprot       ),
      .s_axi4_awvalid ( s_axi_spi_awvalid      ),
      .s_axi4_awready ( s_axi_spi_awready      ),
      .s_axi4_wdata   ( s_axi_spi_wdata        ),
      .s_axi4_wstrb   ( s_axi_spi_wstrb        ),
      .s_axi4_wlast   ( s_axi_spi_wlast        ),
      .s_axi4_wvalid  ( s_axi_spi_wvalid       ),
      .s_axi4_wready  ( s_axi_spi_wready       ),
      .s_axi4_bresp   ( s_axi_spi_bresp        ),
      .s_axi4_bvalid  ( s_axi_spi_bvalid       ),
      .s_axi4_bready  ( s_axi_spi_bready       ),
      .s_axi4_araddr  ( s_axi_spi_araddr[23:0] ),
      .s_axi4_arlen   ( s_axi_spi_arlen        ),
      .s_axi4_arsize  ( s_axi_spi_arsize       ),
      .s_axi4_arburst ( s_axi_spi_arburst      ),
      .s_axi4_arlock  ( s_axi_spi_arlock       ),
      .s_axi4_arcache ( s_axi_spi_arcache      ),
      .s_axi4_arprot  ( s_axi_spi_arprot       ),
      .s_axi4_arvalid ( s_axi_spi_arvalid      ),
      .s_axi4_arready ( s_axi_spi_arready      ),
      .s_axi4_rdata   ( s_axi_spi_rdata        ),
      .s_axi4_rresp   ( s_axi_spi_rresp        ),
      .s_axi4_rlast   ( s_axi_spi_rlast        ),
      .s_axi4_rvalid  ( s_axi_spi_rvalid       ),
      .s_axi4_rready  ( s_axi_spi_rready       ),
      .io0_i          ( '0                     ),
      .io0_o          ( spi_mosi               ),
      .io0_t          (                        ),
      .io1_i          ( spi_miso               ),
      .io1_o          (                        ),
      .io1_t          (                        ),
      .ss_i           ( '0                     ),
      .ss_o           ( spi_ss                 ),
      .ss_t           (                        ),
      .sck_o          ( spi_clk_o              ),
      .sck_i          ( '0                     ),
      .sck_t          (                        ),
      .ip2intc_irpt   ( irq_sources[1]         )
    );
  end else begin
    assign spi_clk_o = 1'b0;
    assign spi_mosi = 1'b0;
    assign spi_ss = 1'b0;

    // assign irq_sources [1] = 1'b0;
    assign spi.aw_ready = 1'b1;
    assign spi.ar_ready = 1'b1;
    assign spi.w_ready = 1'b1;

    assign spi.b_valid = spi.aw_valid;
    assign spi.b_id = spi.aw_id;
    assign spi.b_resp = axi_pkg::RESP_SLVERR;
    assign spi.b_user = '0;

    assign spi.r_valid = spi.ar_valid;
    assign spi.r_resp = axi_pkg::RESP_SLVERR;
    assign spi.r_data = 'hdeadbeef;
    assign spi.r_last = 1'b1;
  end


  // ---------------
  // 4. Ethernet
  // ---------------
  if (InclEthernet) begin : gen_ethernet

    logic                       clk_200_int, clk_rgmii, clk_rgmii_quad;
    logic                       eth_en, eth_we, eth_int_n, eth_pme_n, eth_mdio_i, eth_mdio_o, eth_mdio_oe;
    logic [AxiAddrWidth-1:0]    eth_addr;
    logic [AxiDataWidth-1:0]    eth_wrdata, eth_rdata;
    logic [AxiDataWidth/8-1:0]  eth_be;

    axi2mem #(
      .AXI_ID_WIDTH   ( AxiIdWidth      ),
      .AXI_ADDR_WIDTH ( AxiAddrWidth    ),
      .AXI_DATA_WIDTH ( AxiDataWidth    ),
      .AXI_USER_WIDTH ( AxiUserWidth    )
    ) i_axi2rom (
      .clk_i  ( clk_i                   ),
      .rst_ni ( rst_ni                  ),
      .slave  ( ethernet                ),
      .req_o  ( eth_en                  ),
      .we_o   ( eth_we                  ),
      .addr_o ( eth_addr                ),
      .be_o   ( eth_be                  ),
      .data_o ( eth_wrdata              ),
      .data_i ( eth_rdata               )
    );

    framing_top eth_rgmii (
      .msoc_clk(clk_i),
      .core_lsu_addr(eth_addr[14:0]),
      .core_lsu_wdata(eth_wrdata),
      .core_lsu_be(eth_be),
      .ce_d(eth_en),
      .we_d(eth_en & eth_we),
      .framing_sel(eth_en),
      .framing_rdata(eth_rdata),
      .rst_int(!rst_ni),
      .clk_int(phy_tx_clk_i), // 125 MHz in-phase
      .clk90_int(eth_clk_i),    // 125 MHz quadrature
      .clk_200_int(clk_200MHz_i),
      /*
      * Ethernet: 1000BASE-T RGMII
      */
      .phy_rx_clk(eth_rxck),
      .phy_rxd(eth_rxd),
      .phy_rx_ctl(eth_rxctl),
      .phy_tx_clk(eth_txck),
      .phy_txd(eth_txd),
      .phy_tx_ctl(eth_txctl),
      .phy_reset_n(eth_rst_n),
      .phy_int_n(eth_int_n),
      .phy_pme_n(eth_pme_n),
      .phy_mdc(eth_mdc),
      .phy_mdio_i(eth_mdio_i),
      .phy_mdio_o(eth_mdio_o),
      .phy_mdio_oe(eth_mdio_oe),
      .eth_irq(irq_sources[2])
    );

    IOBUF #(
      .DRIVE(12), // Specify the output drive strength
      .IBUF_LOW_PWR("TRUE"),  // Low Power - "TRUE", High Performance = "FALSE"
      .IOSTANDARD("DEFAULT"), // Specify the I/O standard
      .SLEW("SLOW") // Specify the output slew rate
    ) IOBUF_inst (
      .O(eth_mdio_i),     // Buffer output
      .IO(eth_mdio),   // Buffer inout port (connect directly to top-level port)
      .I(eth_mdio_o),     // Buffer input
      .T(~eth_mdio_oe)      // 3-state enable input, high=input, low=output
    );

  end else begin
    assign irq_sources [2] = 1'b0;
    assign ethernet.aw_ready = 1'b1;
    assign ethernet.ar_ready = 1'b1;
    assign ethernet.w_ready = 1'b1;

    assign ethernet.b_valid = ethernet.aw_valid;
    assign ethernet.b_id = ethernet.aw_id;
    assign ethernet.b_resp = axi_pkg::RESP_SLVERR;
    assign ethernet.b_user = '0;

    assign ethernet.r_valid = ethernet.ar_valid;
    assign ethernet.r_resp = axi_pkg::RESP_SLVERR;
    assign ethernet.r_data = 'hdeadbeef;
    assign ethernet.r_last = 1'b1;
  end

  // ---------------
  // 5. GPIO 
  // ---------------
  assign gpio.b_user = 1'b0;
  assign gpio.r_user = 1'b0;

  if (InclGPIO) begin : gen_gpio

    logic [31:0] s_axi_gpio_awaddr;
    logic [7:0]  s_axi_gpio_awlen;
    logic [2:0]  s_axi_gpio_awsize;
    logic [1:0]  s_axi_gpio_awburst;
    logic [3:0]  s_axi_gpio_awcache;
    logic        s_axi_gpio_awvalid;
    logic        s_axi_gpio_awready;
    logic [31:0] s_axi_gpio_wdata;
    logic [3:0]  s_axi_gpio_wstrb;
    logic        s_axi_gpio_wvalid;
    logic        s_axi_gpio_wready;
    logic [1:0]  s_axi_gpio_bresp;
    logic        s_axi_gpio_bvalid;
    logic        s_axi_gpio_bready;
    logic [31:0] s_axi_gpio_araddr;
    logic [7:0]  s_axi_gpio_arlen;
    logic [2:0]  s_axi_gpio_arsize;
    logic [1:0]  s_axi_gpio_arburst;
    logic [3:0]  s_axi_gpio_arcache;
    logic        s_axi_gpio_arvalid;
    logic        s_axi_gpio_arready;
    logic [31:0] s_axi_gpio_rdata;
    logic [1:0]  s_axi_gpio_rresp;
    logic        s_axi_gpio_rlast;
    logic        s_axi_gpio_rvalid;
    logic        s_axi_gpio_rready;

    // system-bus is 64-bit, convert down to 32 bit
    xlnx_axi_dwidth_converter i_xlnx_axi_dwidth_converter_gpio (
      .s_axi_aclk     ( clk_i              ),
      .s_axi_aresetn  ( rst_ni             ),
      .s_axi_awid     ( gpio.aw_id         ),
      .s_axi_awaddr   ( gpio.aw_addr[31:0] ),
      .s_axi_awlen    ( gpio.aw_len        ),
      .s_axi_awsize   ( gpio.aw_size       ),
      .s_axi_awburst  ( gpio.aw_burst      ),
      .s_axi_awlock   ( gpio.aw_lock       ),
      .s_axi_awcache  ( gpio.aw_cache      ),
      .s_axi_awprot   ( gpio.aw_prot       ),
      .s_axi_awregion ( gpio.aw_region     ),
      .s_axi_awqos    ( gpio.aw_qos        ),
      .s_axi_awvalid  ( gpio.aw_valid      ),
      .s_axi_awready  ( gpio.aw_ready      ),
      .s_axi_wdata    ( gpio.w_data        ),
      .s_axi_wstrb    ( gpio.w_strb        ),
      .s_axi_wlast    ( gpio.w_last        ),
      .s_axi_wvalid   ( gpio.w_valid       ),
      .s_axi_wready   ( gpio.w_ready       ),
      .s_axi_bid      ( gpio.b_id          ),
      .s_axi_bresp    ( gpio.b_resp        ),
      .s_axi_bvalid   ( gpio.b_valid       ),
      .s_axi_bready   ( gpio.b_ready       ),
      .s_axi_arid     ( gpio.ar_id         ),
      .s_axi_araddr   ( gpio.ar_addr[31:0] ),
      .s_axi_arlen    ( gpio.ar_len        ),
      .s_axi_arsize   ( gpio.ar_size       ),
      .s_axi_arburst  ( gpio.ar_burst      ),
      .s_axi_arlock   ( gpio.ar_lock       ),
      .s_axi_arcache  ( gpio.ar_cache      ),
      .s_axi_arprot   ( gpio.ar_prot       ),
      .s_axi_arregion ( gpio.ar_region     ),
      .s_axi_arqos    ( gpio.ar_qos        ),
      .s_axi_arvalid  ( gpio.ar_valid      ),
      .s_axi_arready  ( gpio.ar_ready      ),
      .s_axi_rid      ( gpio.r_id          ),
      .s_axi_rdata    ( gpio.r_data        ),
      .s_axi_rresp    ( gpio.r_resp        ),
      .s_axi_rlast    ( gpio.r_last        ),
      .s_axi_rvalid   ( gpio.r_valid       ),
      .s_axi_rready   ( gpio.r_ready       ),

      .m_axi_awaddr   ( s_axi_gpio_awaddr  ),
      .m_axi_awlen    ( s_axi_gpio_awlen   ),
      .m_axi_awsize   ( s_axi_gpio_awsize  ),
      .m_axi_awburst  ( s_axi_gpio_awburst ),
      .m_axi_awlock   (                    ),
      .m_axi_awcache  ( s_axi_gpio_awcache ),
      .m_axi_awprot   (                    ),
      .m_axi_awregion (                    ),
      .m_axi_awqos    (                    ),
      .m_axi_awvalid  ( s_axi_gpio_awvalid ),
      .m_axi_awready  ( s_axi_gpio_awready ),
      .m_axi_wdata    ( s_axi_gpio_wdata   ),
      .m_axi_wstrb    ( s_axi_gpio_wstrb   ),
      .m_axi_wlast    (                    ),
      .m_axi_wvalid   ( s_axi_gpio_wvalid  ),
      .m_axi_wready   ( s_axi_gpio_wready  ),
      .m_axi_bresp    ( s_axi_gpio_bresp   ),
      .m_axi_bvalid   ( s_axi_gpio_bvalid  ),
      .m_axi_bready   ( s_axi_gpio_bready  ),
      .m_axi_araddr   ( s_axi_gpio_araddr  ),
      .m_axi_arlen    ( s_axi_gpio_arlen   ),
      .m_axi_arsize   ( s_axi_gpio_arsize  ),
      .m_axi_arburst  ( s_axi_gpio_arburst ),
      .m_axi_arlock   (                    ),
      .m_axi_arcache  ( s_axi_gpio_arcache ),
      .m_axi_arprot   (                    ),
      .m_axi_arregion (                    ),
      .m_axi_arqos    (                    ),
      .m_axi_arvalid  ( s_axi_gpio_arvalid ),
      .m_axi_arready  ( s_axi_gpio_arready ),
      .m_axi_rdata    ( s_axi_gpio_rdata   ),
      .m_axi_rresp    ( s_axi_gpio_rresp   ),
      .m_axi_rlast    ( s_axi_gpio_rlast   ),
      .m_axi_rvalid   ( s_axi_gpio_rvalid  ),
      .m_axi_rready   ( s_axi_gpio_rready  )
    );

    xlnx_axi_gpio i_xlnx_axi_gpio (
      .s_axi_aclk    ( clk_i                  ),
      .s_axi_aresetn ( rst_ni                 ),
      .s_axi_awaddr  ( s_axi_gpio_awaddr[8:0] ),
      .s_axi_awvalid ( s_axi_gpio_awvalid     ),
      .s_axi_awready ( s_axi_gpio_awready     ),
      .s_axi_wdata   ( s_axi_gpio_wdata       ),
      .s_axi_wstrb   ( s_axi_gpio_wstrb       ),
      .s_axi_wvalid  ( s_axi_gpio_wvalid      ),
      .s_axi_wready  ( s_axi_gpio_wready      ),
      .s_axi_bresp   ( s_axi_gpio_bresp       ),
      .s_axi_bvalid  ( s_axi_gpio_bvalid      ),
      .s_axi_bready  ( s_axi_gpio_bready      ),
      .s_axi_araddr  ( s_axi_gpio_araddr[8:0] ),
      .s_axi_arvalid ( s_axi_gpio_arvalid     ),
      .s_axi_arready ( s_axi_gpio_arready     ),
      .s_axi_rdata   ( s_axi_gpio_rdata       ),
      .s_axi_rresp   ( s_axi_gpio_rresp       ),
      .s_axi_rvalid  ( s_axi_gpio_rvalid      ),
      .s_axi_rready  ( s_axi_gpio_rready      ),
      .gpio_io_i     ( '0                     ),
      .gpio_io_o     ( leds_o                 ),
      .gpio_io_t     (                        ),
      .gpio2_io_i    ( dip_switches_i         )
    );

    assign s_axi_gpio_rlast = 1'b1;

  end

  // ---------------
  // 6. Timer 
  // ---------------
  if (InclTimer) begin : gen_timer
    logic         timer_penable;
    logic         timer_pwrite;
    logic [31:0]  timer_paddr;
    logic         timer_psel;
    logic [31:0]  timer_pwdata;
    logic [31:0]  timer_prdata;
    logic         timer_pready;
    logic         timer_pslverr;

    axi2apb_64_32 #(
      .AXI4_ADDRESS_WIDTH ( AxiAddrWidth ),
      .AXI4_RDATA_WIDTH   ( AxiDataWidth ),
      .AXI4_WDATA_WIDTH   ( AxiDataWidth ),
      .AXI4_ID_WIDTH      ( AxiIdWidth   ),
      .AXI4_USER_WIDTH    ( AxiUserWidth ),
      .BUFF_DEPTH_SLAVE   ( 2            ),
      .APB_ADDR_WIDTH     ( 32           )
    ) i_axi2apb_64_32_timer (
      .ACLK      ( clk_i           ),
      .ARESETn   ( rst_ni          ),
      .test_en_i ( 1'b0            ),
      .AWID_i    ( timer.aw_id     ),
      .AWADDR_i  ( timer.aw_addr   ),
      .AWLEN_i   ( timer.aw_len    ),
      .AWSIZE_i  ( timer.aw_size   ),
      .AWBURST_i ( timer.aw_burst  ),
      .AWLOCK_i  ( timer.aw_lock   ),
      .AWCACHE_i ( timer.aw_cache  ),
      .AWPROT_i  ( timer.aw_prot   ),
      .AWREGION_i( timer.aw_region ),
      .AWUSER_i  ( timer.aw_user   ),
      .AWQOS_i   ( timer.aw_qos    ),
      .AWVALID_i ( timer.aw_valid  ),
      .AWREADY_o ( timer.aw_ready  ),
      .WDATA_i   ( timer.w_data    ),
      .WSTRB_i   ( timer.w_strb    ),
      .WLAST_i   ( timer.w_last    ),
      .WUSER_i   ( timer.w_user    ),
      .WVALID_i  ( timer.w_valid   ),
      .WREADY_o  ( timer.w_ready   ),
      .BID_o     ( timer.b_id      ),
      .BRESP_o   ( timer.b_resp    ),
      .BVALID_o  ( timer.b_valid   ),
      .BUSER_o   ( timer.b_user    ),
      .BREADY_i  ( timer.b_ready   ),
      .ARID_i    ( timer.ar_id     ),
      .ARADDR_i  ( timer.ar_addr   ),
      .ARLEN_i   ( timer.ar_len    ),
      .ARSIZE_i  ( timer.ar_size   ),
      .ARBURST_i ( timer.ar_burst  ),
      .ARLOCK_i  ( timer.ar_lock   ),
      .ARCACHE_i ( timer.ar_cache  ),
      .ARPROT_i  ( timer.ar_prot   ),
      .ARREGION_i( timer.ar_region ),
      .ARUSER_i  ( timer.ar_user   ),
      .ARQOS_i   ( timer.ar_qos    ),
      .ARVALID_i ( timer.ar_valid  ),
      .ARREADY_o ( timer.ar_ready  ),
      .RID_o     ( timer.r_id      ),
      .RDATA_o   ( timer.r_data    ),
      .RRESP_o   ( timer.r_resp    ),
      .RLAST_o   ( timer.r_last    ),
      .RUSER_o   ( timer.r_user    ),
      .RVALID_o  ( timer.r_valid   ),
      .RREADY_i  ( timer.r_ready   ),
      .PENABLE   ( timer_penable   ),
      .PWRITE    ( timer_pwrite    ),
      .PADDR     ( timer_paddr     ),
      .PSEL      ( timer_psel      ),
      .PWDATA    ( timer_pwdata    ),
      .PRDATA    ( timer_prdata    ),
      .PREADY    ( timer_pready    ),
      .PSLVERR   ( timer_pslverr   )
    );

    apb_timer #(
      .APB_ADDR_WIDTH ( 32 ),
      .TIMER_CNT      ( 2  )
    ) i_timer (
      .HCLK    ( clk_i            ),
      .HRESETn ( rst_ni           ),
      .PSEL    ( timer_psel       ),
      .PENABLE ( timer_penable    ),
      .PWRITE  ( timer_pwrite     ),
      .PADDR   ( timer_paddr      ),
      .PWDATA  ( timer_pwdata     ),
      .PRDATA  ( timer_prdata     ),
      .PREADY  ( timer_pready     ),
      .PSLVERR ( timer_pslverr    ),
      .irq_o   ( irq_sources[6:3] )
    );
  end

  // ---------------
  // 7. VGA 
  // ---------------

  // RegBus interface
    
  // RegBus parameters
  localparam int unsigned RegBusAddrWidth = 32;
  localparam int unsigned RegBusDataWidth = 32;
  localparam int unsigned RegBusStrbWidth =  4;
  localparam int unsigned AXIStrbWidth  =  8;
  
  
  `REG_BUS_TYPEDEF_ALL(reg_vga, logic [RegBusAddrWidth-1:0], logic [RegBusDataWidth-1:0], logic [RegBusStrbWidth-1:0])
  
  REG_BUS #(
    .ADDR_WIDTH ( RegBusAddrWidth  ),
    .DATA_WIDTH ( RegBusDataWidth  )
  ) i_vga_regbus (clk_i );

  reg_vga_req_t vga_reg_req;
  reg_vga_rsp_t vga_reg_rsp;
  
  `REG_BUS_ASSIGN_TO_REQ(vga_reg_req, i_vga_regbus)
  `REG_BUS_ASSIGN_FROM_RSP(i_vga_regbus, vga_reg_rsp)
   
  logic         vga_penable;
  logic         vga_pwrite;
  logic [31:0]  vga_paddr;
  logic         vga_psel;
  logic [31:0]  vga_pwdata;
  logic [31:0]  vga_prdata;
  logic         vga_pready;
  logic         vga_pslverr;

  axi2apb_64_32 #(
    .AXI4_ADDRESS_WIDTH ( AxiAddrWidth  ),
    .AXI4_RDATA_WIDTH   ( AxiDataWidth  ),
    .AXI4_WDATA_WIDTH   ( AxiDataWidth  ),
    .AXI4_ID_WIDTH      ( AxiIdWidth    ),
    .AXI4_USER_WIDTH    ( AxiUserWidth  ),
    .BUFF_DEPTH_SLAVE   ( 2             ),
    .APB_ADDR_WIDTH     ( 32            )
  ) i_axi2apb_64_32_vga (
    .ACLK      ( clk_i          ),
    .ARESETn   ( rst_ni         ),
    .test_en_i ( 1'b0           ),
    .AWID_i    ( vga.aw_id     ),
    .AWADDR_i  ( vga.aw_addr   ),
    .AWLEN_i   ( vga.aw_len    ),
    .AWSIZE_i  ( vga.aw_size   ),
    .AWBURST_i ( vga.aw_burst  ),
    .AWLOCK_i  ( vga.aw_lock   ),
    .AWCACHE_i ( vga.aw_cache  ),
    .AWPROT_i  ( vga.aw_prot   ),
    .AWREGION_i( vga.aw_region ),
    .AWUSER_i  ( vga.aw_user   ),
    .AWQOS_i   ( vga.aw_qos    ),
    .AWVALID_i ( vga.aw_valid  ),
    .AWREADY_o ( vga.aw_ready  ),
    .WDATA_i   ( vga.w_data    ),
    .WSTRB_i   ( vga.w_strb    ),
    .WLAST_i   ( vga.w_last    ),
    .WUSER_i   ( vga.w_user    ),
    .WVALID_i  ( vga.w_valid   ),
    .WREADY_o  ( vga.w_ready   ),
    .BID_o     ( vga.b_id      ),
    .BRESP_o   ( vga.b_resp    ),
    .BVALID_o  ( vga.b_valid   ),
    .BUSER_o   ( vga.b_user    ),
    .BREADY_i  ( vga.b_ready   ),
    .ARID_i    ( vga.ar_id     ),
    .ARADDR_i  ( vga.ar_addr   ),
    .ARLEN_i   ( vga.ar_len    ),
    .ARSIZE_i  ( vga.ar_size   ),
    .ARBURST_i ( vga.ar_burst  ),
    .ARLOCK_i  ( vga.ar_lock   ),
    .ARCACHE_i ( vga.ar_cache  ),
    .ARPROT_i  ( vga.ar_prot   ),
    .ARREGION_i( vga.ar_region ),
    .ARUSER_i  ( vga.ar_user   ),
    .ARQOS_i   ( vga.ar_qos    ),
    .ARVALID_i ( vga.ar_valid  ),
    .ARREADY_o ( vga.ar_ready  ),
    .RID_o     ( vga.r_id      ),
    .RDATA_o   ( vga.r_data    ),
    .RRESP_o   ( vga.r_resp    ),
    .RLAST_o   ( vga.r_last    ),
    .RUSER_o   ( vga.r_user    ),
    .RVALID_o  ( vga.r_valid   ),
    .RREADY_i  ( vga.r_ready   ),
    .PENABLE   ( vga_penable   ),
    .PWRITE    ( vga_pwrite    ),
    .PADDR     ( vga_paddr     ),
    .PSEL      ( vga_psel      ),
    .PWDATA    ( vga_pwdata    ),
    .PRDATA    ( vga_prdata    ),
    .PREADY    ( vga_pready    ),
    .PSLVERR   ( vga_pslverr   )
  );

  apb_to_reg i_apb_to_reg_vga (
    .clk_i     ( clk_i       ),
    .rst_ni    ( rst_ni      ),
    .penable_i ( vga_penable ),
    .pwrite_i  ( vga_pwrite  ),
    .paddr_i   ( vga_paddr   ),
    .psel_i    ( vga_psel    ),
    .pwdata_i  ( vga_pwdata  ),
    .prdata_o  ( vga_prdata  ),
    .pready_o  ( vga_pready  ),
    .pslverr_o ( vga_pslverr ),
    .reg_o     ( i_vga_regbus)
  );
    
  // AXI interface master
  ariane_axi_soc::req_t  vga_axi_req;
  ariane_axi_soc::resp_t vga_axi_resp;
  `AXI_ASSIGN_FROM_REQ(mvga, vga_axi_req)
  `AXI_ASSIGN_TO_RESP(vga_axi_resp, mvga)
    
  // VGA interface
  axi_vga #(
    .RedWidth(   RedWidth)   ,
    .GreenWidth(GreenWidth)    ,
    .BlueWidth(BlueWidth)     ,
    .HCountWidth(HCountWidth)   ,
    .VCountWidth(VCountWidth)   ,
    .AXIAddrWidth   (AxiAddrWidth           ),
    .AXIDataWidth   (AxiDataWidth           ),
    .AXIStrbWidth   (AXIStrbWidth           ),
    .axi_req_t      (ariane_axi_soc::req_t  ),
    .axi_resp_t     (ariane_axi_soc::resp_t ),
    .reg_req_t      (reg_vga_req_t          ),
    .reg_rsp_t      (reg_vga_rsp_t          )
  ) i_axi_vga (
    .clk_i          (clk_i          ),
    .pxl_clk        (clk_vga_i      ),
    .rst_ni         (rst_ni         ),

    .test_mode_en_i (1'b1           ),

    // Regbus config ports
    .reg_req_i      (vga_reg_req   ),
    .reg_rsp_o      (vga_reg_rsp   ),

    // AXI Data ports
    .axi_req_o      (vga_axi_req   ),
    .axi_resp_i     (vga_axi_resp  ),

    // VGA interface
    .hsync_o        (hsync         ),
    .vsync_o        (vsync         ),
    .red_o          (red           ),
    .green_o        (green         ),
    .blue_o         (blue          )
  );

endmodule
