/* Copyright 2018 ETH Zurich and University of Bologna.
 * Copyright and related rights are licensed under the Solderpad Hardware
 * License, Version 0.51 (the "License"); you may not use this file except in
 * compliance with the License.  You may obtain a copy of the License at
 * http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
 * or agreed to in writing, software, hardware and materials distributed under
 * this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
 * CONDITIONS OF ANY KIND, either express or implied. See the License for the
 * specific language governing permissions and limitations under the License.
 *
 * File: $filename.v
 *
 * Description: Auto-generated bootrom
 */

// Auto-generated code
module bootrom_32 (
   input  logic         clk_i,
   input  logic         req_i,
   input  logic [63:0]  addr_i,
   output logic [63:0]  rdata_o
);
    localparam int RomSize = 928;

    const logic [RomSize-1:0][63:0] mem = {
        64'h00000000_0a0d2165,
        64'h6e6f6420_00206567,
        64'h616d6920_746f6f62,
        64'h20676e69_79706f63,
        64'h00000009_3a656d61,
        64'h6e090a0d_00093a73,
        64'h65747562_69727474,
        64'h61090a0d_00000009,
        64'h3a61626c_20747361,
        64'h6c090a0d_0000093a,
        64'h61626c20_74737269,
        64'h66090a0d_00000000,
        64'h09202020_20203a64,
        64'h69756720_6e6f6974,
        64'h69747261_70090a0d,
        64'h00000000_093a6469,
        64'h75672065_70797420,
        64'h6e6f6974_69747261,
        64'h70090a0d_00000000,
        64'h20797274_6e65206e,
        64'h6f697469_74726170,
        64'h20747067_00000009,
        64'h20203a73_65697274,
        64'h6e65206e_6f697469,
        64'h74726170_20657a69,
        64'h73090a0d_00000009,
        64'h3a736569_72746e65,
        64'h206e6f69_74697472,
        64'h61702072_65626d75,
        64'h6e090a0d_00000009,
        64'h2020203a_61626c20,
        64'h73656972_746e6520,
        64'h6e6f6974_69747261,
        64'h70090a0d_00093a61,
        64'h646c2070_756b6361,
        64'h62090a0d_00000000,
        64'h093a6162_6c20746e,
        64'h65727275_63090a0d,
        64'h00000009_3a646576,
        64'h72657365_72090a0d,
        64'h00093a72_65646165,
        64'h685f6372_63090a0d,
        64'h00000909_3a657a69,
        64'h73090a0d_00000009,
        64'h3a6e6f69_73697665,
        64'h72090a0d_0000093a,
        64'h65727574_616e6769,
        64'h73090a0d_003a7265,
        64'h64616568_20656c62,
        64'h6174206e_6f697469,
        64'h74726170_20747067,
        64'h0000203a_65756c61,
        64'h76206e72_75746572,
        64'h2079706f_63206473,
        64'h0000000a_0d216465,
        64'h6c696166_20647261,
        64'h63204453_0000000a,
        64'h0d216465_7a696c61,
        64'h6974696e_69206473,
        64'h00000000_0a0d676e,
        64'h69746978_65202e2e,
        64'h2e647320_657a696c,
        64'h61697469_6e692074,
        64'h6f6e2064_6c756f63,
        64'h0000002e_0000000a,
        64'h0d6b636f_6c622044,
        64'h53206461_65722074,
        64'h6f6e2064_6c756f63,
        64'h0000000a_0d202e2e,
        64'h2e445320_676e697a,
        64'h696c6169_74696e69,
        64'h00000031_34646d63,
        64'h00000035_35646d63,
        64'h00000000_30646d63,
        64'h00000020_3a206573,
        64'h6e6f7073_65720920,
        64'h0020646e_616d6d6f,
        64'h63204453_00000000,
        64'h203f3f79_74706d65,
        64'h20746f6e_206f6669,
        64'h66207872_00000a0d,
        64'h2164657a_696c6169,
        64'h74696e69_20495053,
        64'h00000a0d_00007830,
        64'h203a7375_74617473,
        64'h00000a0d_49505320,
        64'h74696e69_00000a0d,
        64'h21646c72_6f57206f,
        64'h6c6c6548_00000068,
        64'h74646977_2d6f692d,
        64'h67657200_74666968,
        64'h732d6765_72007374,
        64'h70757272_65746e69,
        64'h00746e65_7261702d,
        64'h74707572_7265746e,
        64'h69006465_6570732d,
        64'h746e6572_72756300,
        64'h7665646e_2c766373,
        64'h69720079_7469726f,
        64'h6972702d_78616d2c,
        64'h76637369_72007365,
        64'h6d616e2d_67657200,
        64'h6465646e_65747865,
        64'h2d737470_75727265,
        64'h746e6900_6e6f6967,
        64'h65722d79_726f6d65,
        64'h6d007461_6d726f66,
        64'h0065646f_6d5f6167,
        64'h76006564_69727473,
        64'h00746867_69656800,
        64'h68746469_77006874,
        64'h61702d74_756f6474,
        64'h73007061_6d2d6f6e,
        64'h00736567_6e617200,
        64'h656c646e_61687000,
        64'h72656c6c_6f72746e,
        64'h6f632d74_70757272,
        64'h65746e69_00736c6c,
        64'h65632d74_70757272,
        64'h65746e69_23007469,
        64'h6c70732d_626c7400,
        64'h65707974_2d756d6d,
        64'h00617369_2c766373,
        64'h69720073_75746174,
        64'h73006765_72006570,
        64'h79745f65_63697665,
        64'h64007963_6e657571,
        64'h6572662d_6b636f6c,
        64'h63007963_6e657571,
        64'h6572662d_65736162,
        64'h656d6974_006c6564,
        64'h6f6d0065_6c626974,
        64'h61706d6f_6300736c,
        64'h6c65632d_657a6973,
        64'h2300736c_6c65632d,
        64'h73736572_64646123,
        64'h09000000_02000000,
        64'h02000000_02000000,
        64'h006c6f72_746e6f63,
        64'h11010000_08000000,
        64'h03000000_03000000,
        64'h47010000_04000000,
        64'h03000000_00100000,
        64'h00000018_5b000000,
        64'h08000000_03000000,
        64'h07000000_06000000,
        64'h05000000_04000000,
        64'h58010000_10000000,
        64'h03000000_00007265,
        64'h6d69745f_6270612c,
        64'h706c7570_1b000000,
        64'h0f000000_03000000,
        64'h00003030_30303030,
        64'h38314072_656d6974,
        64'h01000000_02000000,
        64'h04000000_6d010000,
        64'h04000000_03000000,
        64'h02000000_63010000,
        64'h04000000_03000000,
        64'h01000000_58010000,
        64'h04000000_03000000,
        64'h03000000_47010000,
        64'h04000000_03000000,
        64'h00c20100_39010000,
        64'h04000000_03000000,
        64'h80f0fa02_3f000000,
        64'h04000000_03000000,
        64'h00100000_00000010,
        64'h5b000000_08000000,
        64'h03000000_00000000,
        64'h61303535_3631736e,
        64'h1b000000_09000000,
        64'h03000000_00000030,
        64'h30303030_30303140,
        64'h74726175_01000000,
        64'h02000000_03000000,
        64'ha9000000_04000000,
        64'h03000000_1e000000,
        64'h2e010000_04000000,
        64'h03000000_07000000,
        64'h1b010000_04000000,
        64'h03000000_00000004,
        64'h0000000c_5b000000,
        64'h08000000_03000000,
        64'h09000000_02000000,
        64'h0b000000_02000000,
        64'hfd000000_10000000,
        64'h03000000_94000000,
        64'h00000000_03000000,
        64'h00306369_6c702c76,
        64'h63736972_1b000000,
        64'h0c000000_03000000,
        64'h01000000_83000000,
        64'h04000000_03000000,
        64'h00000000_00000000,
        64'h04000000_03000000,
        64'h00000000_30303030,
        64'h30306340_72656c6c,
        64'h6f72746e_6f632d74,
        64'h70757272_65746e69,
        64'h01000000_02000000,
        64'h006c6f72_746e6f63,
        64'h11010000_08000000,
        64'h03000000_00000c00,
        64'h00000002_5b000000,
        64'h08000000_03000000,
        64'h07000000_02000000,
        64'h03000000_02000000,
        64'hfd000000_10000000,
        64'h03000000_00000000,
        64'h30746e69_6c632c76,
        64'h63736972_1b000000,
        64'h0d000000_03000000,
        64'h00000030_30303030,
        64'h30324074_6e696c63,
        64'h01000000_b1000000,
        64'h00000000_03000000,
        64'h00007375_622d656c,
        64'h706d6973_00636f73,
        64'h2d657261_622d656e,
        64'h61697261_2c687465,
        64'h1b000000_1f000000,
        64'h03000000_01000000,
        64'h0f000000_04000000,
        64'h03000000_01000000,
        64'h00000000_04000000,
        64'h03000000_00636f73,
        64'h01000000_02000000,
        64'h02000000_01000000,
        64'hef000000_04000000,
        64'h03000000_80f0fa02,
        64'h3f000000_04000000,
        64'h03000000_00003562,
        64'h36673572_e8000000,
        64'h07000000_03000000,
        64'h00000000_df000000,
        64'h04000000_03000000,
        64'h00050000_d8000000,
        64'h04000000_03000000,
        64'he0010000_d1000000,
        64'h04000000_03000000,
        64'h80020000_cb000000,
        64'h04000000_03000000,
        64'h00100000_00000050,
        64'h00600900_000000a0,
        64'h5b000000_10000000,
        64'h03000000_00000000,
        64'h72656666_7562656d,
        64'h6172662d_61677663,
        64'h1b000000_11000000,
        64'h03000000_00000000,
        64'h30303030_30303061,
        64'h40616776_01000000,
        64'hb1000000_00000000,
        64'h03000000_01000000,
        64'h0f000000_04000000,
        64'h03000000_01000000,
        64'h00000000_04000000,
        64'h03000000_00000030,
        64'h30323531_313a3030,
        64'h30303030_30314074,
        64'h7261752f_636f732f,
        64'hbf000000_1a000000,
        64'h03000000_00006e65,
        64'h736f6863_01000000,
        64'h02000000_02000000,
        64'h01000000_a9000000,
        64'h04000000_03000000,
        64'h00000010_000000a0,
        64'h5b000000_08000000,
        64'h03000000_b8000000,
        64'h00000000_03000000,
        64'h00000000_30407265,
        64'h66667562_01000000,
        64'hb1000000_00000000,
        64'h03000000_01000000,
        64'h0f000000_04000000,
        64'h03000000_01000000,
        64'h00000000_04000000,
        64'h03000000_0079726f,
        64'h6d656d2d_64657672,
        64'h65736572_01000000,
        64'h02000000_00000040,
        64'h00000080_5b000000,
        64'h08000000_03000000,
        64'h00007972_6f6d656d,
        64'h4f000000_07000000,
        64'h03000000_00303030,
        64'h30303030_38407972,
        64'h6f6d656d_01000000,
        64'h02000000_02000000,
        64'h02000000_02000000,
        64'ha9000000_04000000,
        64'h03000000_00006374,
        64'h6e692d75_70632c76,
        64'h63736972_1b000000,
        64'h0f000000_03000000,
        64'h94000000_00000000,
        64'h03000000_01000000,
        64'h83000000_04000000,
        64'h03000000_00000000,
        64'h72656c6c_6f72746e,
        64'h6f632d74_70757272,
        64'h65746e69_01000000,
        64'h79000000_00000000,
        64'h03000000_00003233,
        64'h76732c76_63736972,
        64'h70000000_0b000000,
        64'h03000000_00616d69,
        64'h32337672_66000000,
        64'h08000000_03000000,
        64'h00000076_63736972,
        64'h00656e61_69726120,
        64'h2c687465_1b000000,
        64'h12000000_03000000,
        64'h00000000_79616b6f,
        64'h5f000000_05000000,
        64'h03000000_00000000,
        64'h5b000000_04000000,
        64'h03000000_00757063,
        64'h4f000000_04000000,
        64'h03000000_80f0fa02,
        64'h3f000000_04000000,
        64'h03000000_00000030,
        64'h40757063_01000000,
        64'h40787d01_2c000000,
        64'h04000000_03000000,
        64'h00000000_0f000000,
        64'h04000000_03000000,
        64'h01000000_00000000,
        64'h04000000_03000000,
        64'h00000000_73757063,
        64'h01000000_00657261,
        64'h622d656e_61697261,
        64'h2c687465_26000000,
        64'h10000000_03000000,
        64'h00766564_2d657261,
        64'h622d656e_61697261,
        64'h2c687465_1b000000,
        64'h14000000_03000000,
        64'h01000000_0f000000,
        64'h04000000_03000000,
        64'h01000000_00000000,
        64'h04000000_03000000,
        64'h00000000_01000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h88060000_7a010000,
        64'h00000000_10000000,
        64'h11000000_28000000,
        64'hc0060000_38000000,
        64'h3a080000_edfe0dd0,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h46454443_42413938,
        64'h37363534_33323130,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_0000006f,
        64'h940ff0ef_9e850513,
        64'h00001517_8f4ff0ef,
        64'h00112623_20058593,
        64'h08050513_ff010113,
        64'h02faf537_0001c5b7,
        64'hf11ff06f_ffe00493,
        64'h970ff0ef_a4050513,
        64'h00001517_a44ff0ef,
        64'h41f4d593_00048513,
        64'h988ff0ef_b4450513,
        64'h00001517_994ff0ef,
        64'hb3c50513_00001517,
        64'hf49ff06f_ffe00493,
        64'h9a8ff0ef_a7850513,
        64'h00001517_a7cff0ef,
        64'h41fad593_000a8513,
        64'h9c0ff0ef_b7c50513,
        64'h00001517_9ccff0ef,
        64'hb7450513_00001517,
        64'hf81ff06f_ffe00493,
        64'h9e0ff0ef_ab050513,
        64'h00001517_ab4ff0ef,
        64'h41f4d593_00048513,
        64'h9f8ff0ef_bb450513,
        64'h00001517_a04ff0ef,
        64'hbac50513_00001517,
        64'hfb9ff06f_fff00493,
        64'ha18ff0ef_b8450513,
        64'h00001517_00008067,
        64'h03010113_00812c03,
        64'h00c12b83_01012b03,
        64'h01412a83_01812a03,
        64'h01c12983_02012903,
        64'h02412483_02812403,
        64'h00048513_02c12083,
        64'hfd040113_a5cff0ef,
        64'hdbc50513_00001517,
        64'h04051e63_00050493,
        64'hbb1ff0ef_40b60633,
        64'h00160613_000b8513,
        64'h020c2583_028c2603,
        64'ha88ff0ef_dd450513,
        64'h00001517_f36a94e3,
        64'h080a0a13_08098993,
        64'h08048913_aa4ff0ef,
        64'h001a8a93_b7850513,
        64'h00001517_ff249ae3,
        64'hc0cff0ef_00148493,
        64'h0004c503_ac4ff0ef,
        64'he0450513_00001517,
        64'hb98ff0ef_0149a583,
        64'h0109a503_adcff0ef,
        64'he0c50513_00001517,
        64'hbb0ff0ef_0089a503,
        64'h00c9a583_af4ff0ef,
        64'he1450513_00001517,
        64'hbc8ff0ef_fb890493,
        64'h0009a503_0049a583,
        64'hb10ff0ef_e2050513,
        64'h00001517_ff349ae3,
        64'hc74ff0ef_00148493,
        64'h0004c503_000a0493,
        64'hb30ff0ef_e2450513,
        64'h00001517_ff449ae3,
        64'hc94ff0ef_00148493,
        64'h0004c503_f8090493,
        64'hb50ff0ef_e2850513,
        64'h00001517_cb0ff0ef,
        64'h0ffaf513_b64ff0ef,
        64'he2450513_00001517,
        64'h00400b13_01010a13,
        64'h02010993_08010913,
        64'h1a051663_00050a93,
        64'h00010c13_ccdff0ef,
        64'h00010513_00100613,
        64'he0010113_04892583,
        64'hba0ff0ef_c7050513,
        64'h00001517_c0cff0ef,
        64'h05412503_bb4ff0ef,
        64'he5450513_00001517,
        64'hc20ff0ef_05012503,
        64'hbc8ff0ef_e4850513,
        64'h00001517_c9cff0ef,
        64'h04812503_04c12583,
        64'hbe0ff0ef_e4050513,
        64'h00001517_cb4ff0ef,
        64'h02012503_02412583,
        64'hbf8ff0ef_e4850513,
        64'h00001517_cccff0ef,
        64'h01812503_01c12583,
        64'hc10ff0ef_e4c50513,
        64'h00001517_c7cff0ef,
        64'h01412503_c24ff0ef,
        64'he5050513_00001517,
        64'hc90ff0ef_01012503,
        64'hc38ff0ef_e5450513,
        64'h00001517_ca4ff0ef,
        64'h00c12503_c4cff0ef,
        64'he5c50513_00001517,
        64'hcb8ff0ef_00812503,
        64'hc60ff0ef_e6050513,
        64'h00001517_d34ff0ef,
        64'h00012503_00412583,
        64'hc78ff0ef_e6850513,
        64'h00001517_c84ff0ef,
        64'he5850513_00001517,
        64'h2e051a63_00050493,
        64'h00010913_dddff0ef,
        64'h00010513_00100593,
        64'h00100613_e0010113,
        64'hcb0ff0ef_e4450513,
        64'h00001517_28051e63,
        64'hc81ff0ef_00050b93,
        64'h03010413_01812423,
        64'h01612823_01512a23,
        64'h01412c23_01312e23,
        64'h03212023_02912223,
        64'h02112623_01712623,
        64'h02812423_fd010113,
        64'hfc1ff06f_fff00413,
        64'hd00ff0ef_e4c50513,
        64'h00001517_fe041ae3,
        64'hfa0ff0ef_fff40413,
        64'h0ff00513_00800413,
        64'h00008067_0b010113,
        64'h09412a83_0a012903,
        64'h0a812403_00040513,
        64'h0ac12083_08c12b83,
        64'h09012b03_09812a03,
        64'h09c12983_0a412483,
        64'hfe0ff0ef_0ff00513,
        64'h96dff0ef_00c00513,
        64'h00000593_00100613,
        64'hffe00413_fe5ff06f,
        64'hd70ff0ef_ed850513,
        64'h00001517_0180006f,
        64'h00000413_f32046e3,
        64'hfff90913_00078a63,
        64'h033967b3_03479663,
        64'h000b8a93_0107d793,
        64'h01079793_009567b3,
        64'h839ff0ef_0104d493,
        64'h0ff00513_01049493,
        64'h00851493_84dff0ef,
        64'h0ff00513_f89b94e3,
        64'h040a8a93_040b8b93,
        64'hfada94e3_010a5a13,
        64'h00168693_01079a13,
        64'h00e7c7b3_01677733,
        64'h00579713_4107d793,
        64'h01079793_00e7c7b3,
        64'h00c79713_4107d793,
        64'h01079793_00e7c7b3,
        64'h00f77713_0047d713,
        64'h00e7c7b3_01075713,
        64'h01071713_01476733,
        64'h0006c783_008a5a13,
        64'h008a1713_000b8693,
        64'h981ff0ef_00010513,
        64'h04000593_000b8613,
        64'h200b8493_040a8a93,
        64'h00000a13_000a8b93,
        64'hfe851ce3_8e5ff0ef,
        64'h0ff00513_3e800993,
        64'hfe0b0b13_0fe00413,
        64'h09712623_09412c23,
        64'h0a912223_09312e23,
        64'h00002b37_09612823,
        64'h16051263_a99ff0ef,
        64'h01200513_00100613,
        64'hfed79ce3_00478793,
        64'h00e7a023_fff00713,
        64'h08010693_00010793,
        64'h00060913_00050a93,
        64'h0a812423_0a112623,
        64'h09512a23_0b212023,
        64'hf5010113_00008067,
        64'h01055513_01051513,
        64'h00f54533_00e7f7b3,
        64'hfe070713_00551793,
        64'h00002737_41055513,
        64'h01051513_00f54533,
        64'h00c51793_41055513,
        64'h01051513_00f5c533,
        64'h00f7f793_0045d793,
        64'h00f5c5b3_0107d793,
        64'h01079793_00a7e7b3,
        64'h00855513_00851793,
        64'h00008067_07f57513,
        64'h00f54533_0ff7f793,
        64'h00451793_00b54533,
        64'h00f54533_0045d513,
        64'h0075d793_00b575b3,
        64'hfc1ff06f_ffd00513,
        64'hfc9ff06f_ffe00513,
        64'h00008067_01010113,
        64'hfff00513_00012903,
        64'h00412483_00812403,
        64'h00c12083_00008067,
        64'h01010113_00012903,
        64'h00412483_00812403,
        64'h00c12083_00000513,
        64'h04050263_e7dff0ef,
        64'h04050263_d61ff0ef,
        64'hfa0ff0ef_07050513,
        64'h00001517_901ff0ef,
        64'h00100513_fb4ff0ef,
        64'h0c050513_00001517,
        64'hfc0ff0ef_0dc50513,
        64'h00001517_fccff0ef,
        64'h0cc50513_00001517,
        64'hfd241ee3_06048663,
        64'ha71ff0ef_0ff00513,
        64'hfff48493_00050413,
        64'hc05ff0ef_00000513,
        64'h00000593_09500613,
        64'h00100913_71048493,
        64'h000024b7_fe041ae3,
        64'haa1ff0ef_fff40413,
        64'h0ff00513_00a00413,
        64'h821ff0ef_15450513,
        64'h00001517_9edff0ef,
        64'h01212023_00912223,
        64'h00812423_00112623,
        64'hff010113_00008067,
        64'h01010113_00412483,
        64'h00812403_00143513,
        64'h00c12083_f4940ce3,
        64'haf1ff0ef_0ff00513,
        64'h869ff0ef_13850513,
        64'h00001517_9c9ff0ef,
        64'h00040513_87dff0ef,
        64'h18850513_00001517,
        64'h889ff0ef_1b450513,
        64'h00001517_895ff0ef,
        64'h19450513_00001517,
        64'h00050413_cb9ff0ef,
        64'h02900513_400005b7,
        64'h07700613_8b5ff0ef,
        64'h18450513_00001517,
        64'ha15ff0ef_00040513,
        64'h8c9ff0ef_1d450513,
        64'h00001517_8d5ff0ef,
        64'h1f850513_00001517,
        64'h8e1ff0ef_1e050513,
        64'h00001517_b7dff0ef,
        64'h0ff00513_00050413,
        64'hd0dff0ef_03700513,
        64'h00000593_06500613,
        64'h00100493_00812423,
        64'h00112623_00912223,
        64'hff010113_00008067,
        64'h01010113_00153513,
        64'h00812403_fff40513,
        64'h00c12083_935ff0ef,
        64'h20450513_00001517,
        64'ha95ff0ef_00040513,
        64'h949ff0ef_25450513,
        64'h00001517_955ff0ef,
        64'h27850513_00001517,
        64'h961ff0ef_26050513,
        64'h00001517_bfdff0ef,
        64'h0ff00513_00050413,
        64'hd8dff0ef_00812423,
        64'h00112623_03700513,
        64'h00000593_06500613,
        64'hff010113_00008067,
        64'h01010113_0017b513,
        64'h00012903_00412483,
        64'hf5690793_00812403,
        64'h00c12083_fe8792e3,
        64'h00f4f793_00008067,
        64'h01010113_00012903,
        64'h00412483_00812403,
        64'h00c12083_00f40e63,
        64'h00000513_00100793,
        64'hc71ff0ef_0ff00513,
        64'hc79ff0ef_0ff00513,
        64'h00050913_c85ff0ef,
        64'h0ff00513_00050493,
        64'hc91ff0ef_0ff00513,
        64'hc99ff0ef_0ff00513,
        64'hca1ff0ef_0ff00513,
        64'h00050413_e31ff0ef,
        64'h01212023_00912223,
        64'h00812423_00112623,
        64'h00800513_1aa00593,
        64'h08700613_ff010113,
        64'h00008067_01010113,
        64'h00000513_00012903,
        64'h00412483_00812403,
        64'h00c12083_00008067,
        64'h01010113_00100513,
        64'h00012903_00412483,
        64'h00812403_00c12083,
        64'ha79ff0ef_34850513,
        64'h00001517_bd9ff0ef,
        64'h00100513_a8dff0ef,
        64'h39850513_00001517,
        64'ha99ff0ef_3b450513,
        64'h00001517_aa5ff0ef,
        64'h3a450513_00001517,
        64'hfd241ee3_04048e63,
        64'hd49ff0ef_0ff00513,
        64'hfff48493_00050413,
        64'heddff0ef_00000513,
        64'h00000593_09500613,
        64'h00100913_71048493,
        64'h00812423_00112623,
        64'h01212023_000024b7,
        64'h00912223_ff010113,
        64'haf9ff06f_01010113,
        64'h3cc50513_00001517,
        64'h00412483_00c12083,
        64'h00812403_c69ff0ef,
        64'h00040513_b1dff0ef,
        64'h42850513_00001517,
        64'hb29ff0ef_00048513,
        64'hb31ff0ef_00058413,
        64'h00812423_00112623,
        64'h43c50513_00001517,
        64'h00050493_00912223,
        64'hff010113_00008067,
        64'h01010113_00012903,
        64'h00412483_00812403,
        64'h00c12083_fe07c4e3,
        64'hfff40413_4187d793,
        64'h01851793_e0dff0ef,
        64'h0ff00513_00040e63,
        64'h0080006f_06400413,
        64'he21ff0ef_00048513,
        64'he29ff0ef_0ff47513,
        64'he31ff0ef_0ff57513,
        64'h00845513_e3dff0ef,
        64'h0ff57513_01045513,
        64'he49ff0ef_01845513,
        64'he51ff0ef_04096513,
        64'he59ff0ef_00060493,
        64'h00058413_00912223,
        64'h00812423_00112623,
        64'h0ff00513_00050913,
        64'h01212023_ff010113,
        64'he81ff06f_0ff00513,
        64'h00008067_fff00513,
        64'h00008067_00000513,
        64'h06e7a023_00600713,
        64'h200007b7_06d72823,
        64'hfff00693_20000737,
        64'hfec712e3_feb60fa3,
        64'h00160613_06c7a583,
        64'h200007b7_fe079ae3,
        64'h0017f793_0006a783,
        64'h02c70263_06468693,
        64'h00b60733_200006b7,
        64'hfe079ce3_0017f793,
        64'h00072783_06470713,
        64'h06d7a023_10600693,
        64'h20000737_200007b7,
        64'hfe079ce3_fff78793,
        64'h00000013_03200793,
        64'hfed51ae3_00f72023,
        64'h00150513_00054783,
        64'h00058a63_00b506b3,
        64'h06870713_06d7a823,
        64'h20000737_200007b7,
        64'hffe00693_0ab7e863,
        64'h10000793_fadff06f,
        64'hcb9ff0ef_58850513,
        64'h00001517_d8dff0ef,
        64'h00000593_00042503,
        64'hcd1ff0ef_5b850513,
        64'h00001517_00008067,
        64'h01010113_00412483,
        64'h0ff4f513_06e7a023,
        64'h00600713_200007b7,
        64'h06d72823_fff00693,
        64'h20000737_00812403,
        64'h00c12083_02078a63,
        64'h0017f793_00042783,
        64'h06c72483_20000737,
        64'hfe079ce3_0017f793,
        64'h00042783_06440413,
        64'h06e7a023_10600713,
        64'h20000437_200007b7,
        64'hfe079ce3_fff78793,
        64'h00000013_06a72423,
        64'h06400793_20000737,
        64'h06d7a823_ffe00693,
        64'h200007b7_00912223,
        64'h00812423_00112623,
        64'hff010113_d75ff06f,
        64'h01010113_64c50513,
        64'h00001517_00012903,
        64'h00412483_00c12083,
        64'h00812403_06f42023,
        64'h00600793_d9dff0ef,
        64'h66c50513_00001517,
        64'he71ff0ef_00000593,
        64'h00048513_db5ff0ef,
        64'h67850513_00001517,
        64'h0004a483_06448493,
        64'h06f42023_16600793,
        64'hdd1ff0ef_6a050513,
        64'h00001517_ea5ff0ef,
        64'h00090513_00000593,
        64'hde9ff0ef_6ac50513,
        64'h00001517_0644a903,
        64'h200004b7_06f42023,
        64'h20000437_10400793,
        64'hfe079ce3_fff78793,
        64'h00000013_00a00793,
        64'h04e7a023_00a00713,
        64'h200007b7_e25ff0ef,
        64'h01212023_00912223,
        64'h00812423_00112623,
        64'h6f050513_ff010113,
        64'h00001517_00008067,
        64'h00052503_00008067,
        64'h00b52023_00008067,
        64'h00d78023_100007b7,
        64'hfe078ce3_0207f793,
        64'h00074783_01470713,
        64'h00c78023_100007b7,
        64'h10000737_fe078ce3,
        64'h0207f793_00074783,
        64'h01470713_10000737,
        64'h00074683_0007c603,
        64'h00a787b3_00e78733,
        64'h00455513_00f57713,
        64'he1078793_00001797,
        64'hfa9ff06f_00f6e7b3,
        64'h00c557b3_00df16b3,
        64'h40ce86b3_00008067,
        64'hfbc61ae3_ff860613,
        64'h00688023_fe078ce3,
        64'h0207f793_00074783,
        64'h00d88023_fe078ce3,
        64'h0207f793_00074783,
        64'h0006c683_0007c303,
        64'h00d806b3_00f807b3,
        64'h00f7f793_0046d693,
        64'h0ff7f693_00f5d7b3,
        64'h0407c863_fe060793,
        64'hff800e13_01470713,
        64'h100008b7_01f00e93,
        64'h00159f13_e9c80813,
        64'h03800613_10000737,
        64'h00001817_00008067,
        64'hfa661ee3_ff860613,
        64'h01180023_fe078ce3,
        64'h0207f793_00074783,
        64'h00d80023_fe078ce3,
        64'h0207f793_00074783,
        64'h0006c683_0007c883,
        64'h00d586b3_00f587b3,
        64'h00f7f793_0046d693,
        64'h0ff7f693_00c557b3,
        64'hff800313_01470713,
        64'h10000837_f0458593,
        64'h01800613_10000737,
        64'h00001597_00008067,
        64'h00f58023_0007c783,
        64'h00e580a3_00a787b3,
        64'h00455513_00074703,
        64'h00e78733_00f57713,
        64'hf3078793_00001797,
        64'h00008067_fe0694e3,
        64'h00150513_00154683,
        64'h00d60023_fe078ce3,
        64'h0207f793_00074783,
        64'h01470713_10000637,
        64'h10000737_02068663,
        64'h00054683_00008067,
        64'h00f68823_02000793,
        64'h00f60423_fc700793,
        64'h00e78623_00300713,
        64'h00a70223_0ff57513,
        64'h01058023_00855513,
        64'h0ff57813_100006b7,
        64'h10000637_100005b7,
        64'h00d78623_f8000693,
        64'h100007b7_00070223,
        64'h10000737_02b55533,
        64'h00459593_00008067,
        64'h00a78023_100007b7,
        64'hfe078ce3_0207f793,
        64'h00074783_01470713,
        64'h10000737_00008067,
        64'h02057513_0147c503,
        64'h100007b7_00008067,
        64'h00054503_00008067,
        64'h00b50023_00008067,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00048067_800004b7,
        64'h18858593_00001597,
        64'hf1402573_ff24c6e3,
        64'h40090913_02000937,
        64'h00448493_fe091ee3,
        64'h0004a903_00092023,
        64'h00990933_00291913,
        64'hf1402973_020004b7,
        64'hfe090ae3_00897913,
        64'h34402973_10500073,
        64'hff24c6e3_40090913,
        64'h02000937_00448493,
        64'h0124a023_00100913,
        64'h020004b7_020010ef,
        64'h84000137_03249463,
        64'hf1402973_00000493,
        64'h30491073_00800913
    };

    logic [$clog2(RomSize)-1:0] addr_q;

    always_ff @(posedge clk_i) begin
        if (req_i) begin
            addr_q <= addr_i[$clog2(RomSize)-1+3:3];
        end
    end

    // this prevents spurious Xes from propagating into
    // the speculative fetch stage of the core
    assign rdata_o = (addr_q < RomSize) ? mem[addr_q] : '0;
endmodule
